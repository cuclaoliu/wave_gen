// nios_core.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module nios_core (
		input  wire        altpll_audio_areset_export, // altpll_audio_areset.export
		output wire        altpll_audio_locked_export, // altpll_audio_locked.export
		input  wire        altpll_sys_areset_export,   //   altpll_sys_areset.export
		output wire        altpll_sys_locked_export,   //   altpll_sys_locked.export
		input  wire        audio_bclk,                 //               audio.bclk
		input  wire        audio_adclrc,               //                    .adclrc
		output wire        audio_xck,                  //                    .xck
		input  wire        audio_adcdat,               //                    .adcdat
		input  wire        audio_daclrc,               //                    .daclrc
		output wire        audio_dacdat,               //                    .dacdat
		input  wire        clk_clk,                    //                 clk.clk
		output wire        clk_sdram_clk,              //           clk_sdram.clk
		output wire        clk_vga_clk,                //             clk_vga.clk
		output wire        i2c_scl_export,             //             i2c_scl.export
		inout  wire        i2c_sda_export,             //             i2c_sda.export
		input  wire [3:0]  key_export,                 //                 key.export
		output wire [7:0]  ledg_export,                //                ledg.export
		output wire [15:0] ledr_export,                //                ledr.export
		input  wire        reset_reset_n,              //               reset.reset_n
		input  wire [15:0] sw_export                   //                  sw.export
	);

	wire         altpll_sys_c0_clk;                                         // altpll_sys:c0 -> [clock_crossing_bridge:s0_clk, data_buffer:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:altpll_sys_c0_clk, nios2_gen2:clk, onchip_memory2:clk, rst_controller_003:clk, sysid_qsys:clock, timer:clk]
	wire         altpll_audio_c0_clk;                                       // altpll_audio:c0 -> [audio:clk, mm_interconnect_0:altpll_audio_c0_clk, rst_controller_001:clk]
	wire         altpll_sys_c3_clk;                                         // altpll_sys:c3 -> [clock_crossing_bridge:m0_clk, i2c_scl:clk, i2c_sda:clk, key:clk, ledg:clk, ledr:clk, mm_interconnect_1:altpll_sys_c3_clk, rst_controller_002:clk, sw:clk]
	wire  [31:0] nios2_gen2_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                        // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [24:0] nios2_gen2_data_master_address;                            // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                         // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                               // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire         nios2_gen2_data_master_write;                              // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                          // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [24:0] nios2_gen2_instruction_master_address;                     // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                        // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         nios2_gen2_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [15:0] mm_interconnect_0_audio_avalon_slave_readdata;             // audio:avalon_slave_readdata -> mm_interconnect_0:audio_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_audio_avalon_slave_address;              // mm_interconnect_0:audio_avalon_slave_address -> audio:avalon_slave_address
	wire         mm_interconnect_0_audio_avalon_slave_read;                 // mm_interconnect_0:audio_avalon_slave_read -> audio:avalon_slave_read
	wire         mm_interconnect_0_audio_avalon_slave_write;                // mm_interconnect_0:audio_avalon_slave_write -> audio:avalon_slave_write
	wire  [15:0] mm_interconnect_0_audio_avalon_slave_writedata;            // mm_interconnect_0:audio_avalon_slave_writedata -> audio:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;     // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;  // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_audio_pll_slave_readdata;         // altpll_audio:readdata -> mm_interconnect_0:altpll_audio_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_audio_pll_slave_address;          // mm_interconnect_0:altpll_audio_pll_slave_address -> altpll_audio:address
	wire         mm_interconnect_0_altpll_audio_pll_slave_read;             // mm_interconnect_0:altpll_audio_pll_slave_read -> altpll_audio:read
	wire         mm_interconnect_0_altpll_audio_pll_slave_write;            // mm_interconnect_0:altpll_audio_pll_slave_write -> altpll_audio:write
	wire  [31:0] mm_interconnect_0_altpll_audio_pll_slave_writedata;        // mm_interconnect_0:altpll_audio_pll_slave_writedata -> altpll_audio:writedata
	wire  [31:0] mm_interconnect_0_altpll_sys_pll_slave_readdata;           // altpll_sys:readdata -> mm_interconnect_0:altpll_sys_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_sys_pll_slave_address;            // mm_interconnect_0:altpll_sys_pll_slave_address -> altpll_sys:address
	wire         mm_interconnect_0_altpll_sys_pll_slave_read;               // mm_interconnect_0:altpll_sys_pll_slave_read -> altpll_sys:read
	wire         mm_interconnect_0_altpll_sys_pll_slave_write;              // mm_interconnect_0:altpll_sys_pll_slave_write -> altpll_sys:write
	wire  [31:0] mm_interconnect_0_altpll_sys_pll_slave_writedata;          // mm_interconnect_0:altpll_sys_pll_slave_writedata -> altpll_sys:writedata
	wire  [31:0] mm_interconnect_0_clock_crossing_bridge_s0_readdata;       // clock_crossing_bridge:s0_readdata -> mm_interconnect_0:clock_crossing_bridge_s0_readdata
	wire         mm_interconnect_0_clock_crossing_bridge_s0_waitrequest;    // clock_crossing_bridge:s0_waitrequest -> mm_interconnect_0:clock_crossing_bridge_s0_waitrequest
	wire         mm_interconnect_0_clock_crossing_bridge_s0_debugaccess;    // mm_interconnect_0:clock_crossing_bridge_s0_debugaccess -> clock_crossing_bridge:s0_debugaccess
	wire   [8:0] mm_interconnect_0_clock_crossing_bridge_s0_address;        // mm_interconnect_0:clock_crossing_bridge_s0_address -> clock_crossing_bridge:s0_address
	wire         mm_interconnect_0_clock_crossing_bridge_s0_read;           // mm_interconnect_0:clock_crossing_bridge_s0_read -> clock_crossing_bridge:s0_read
	wire   [3:0] mm_interconnect_0_clock_crossing_bridge_s0_byteenable;     // mm_interconnect_0:clock_crossing_bridge_s0_byteenable -> clock_crossing_bridge:s0_byteenable
	wire         mm_interconnect_0_clock_crossing_bridge_s0_readdatavalid;  // clock_crossing_bridge:s0_readdatavalid -> mm_interconnect_0:clock_crossing_bridge_s0_readdatavalid
	wire         mm_interconnect_0_clock_crossing_bridge_s0_write;          // mm_interconnect_0:clock_crossing_bridge_s0_write -> clock_crossing_bridge:s0_write
	wire  [31:0] mm_interconnect_0_clock_crossing_bridge_s0_writedata;      // mm_interconnect_0:clock_crossing_bridge_s0_writedata -> clock_crossing_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_clock_crossing_bridge_s0_burstcount;     // mm_interconnect_0:clock_crossing_bridge_s0_burstcount -> clock_crossing_bridge:s0_burstcount
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_data_buffer_s1_chipselect;               // mm_interconnect_0:data_buffer_s1_chipselect -> data_buffer:chipselect
	wire  [31:0] mm_interconnect_0_data_buffer_s1_readdata;                 // data_buffer:readdata -> mm_interconnect_0:data_buffer_s1_readdata
	wire   [9:0] mm_interconnect_0_data_buffer_s1_address;                  // mm_interconnect_0:data_buffer_s1_address -> data_buffer:address
	wire   [3:0] mm_interconnect_0_data_buffer_s1_byteenable;               // mm_interconnect_0:data_buffer_s1_byteenable -> data_buffer:byteenable
	wire         mm_interconnect_0_data_buffer_s1_write;                    // mm_interconnect_0:data_buffer_s1_write -> data_buffer:write
	wire  [31:0] mm_interconnect_0_data_buffer_s1_writedata;                // mm_interconnect_0:data_buffer_s1_writedata -> data_buffer:writedata
	wire         mm_interconnect_0_data_buffer_s1_clken;                    // mm_interconnect_0:data_buffer_s1_clken -> data_buffer:clken
	wire         clock_crossing_bridge_m0_waitrequest;                      // mm_interconnect_1:clock_crossing_bridge_m0_waitrequest -> clock_crossing_bridge:m0_waitrequest
	wire  [31:0] clock_crossing_bridge_m0_readdata;                         // mm_interconnect_1:clock_crossing_bridge_m0_readdata -> clock_crossing_bridge:m0_readdata
	wire         clock_crossing_bridge_m0_debugaccess;                      // clock_crossing_bridge:m0_debugaccess -> mm_interconnect_1:clock_crossing_bridge_m0_debugaccess
	wire   [8:0] clock_crossing_bridge_m0_address;                          // clock_crossing_bridge:m0_address -> mm_interconnect_1:clock_crossing_bridge_m0_address
	wire         clock_crossing_bridge_m0_read;                             // clock_crossing_bridge:m0_read -> mm_interconnect_1:clock_crossing_bridge_m0_read
	wire   [3:0] clock_crossing_bridge_m0_byteenable;                       // clock_crossing_bridge:m0_byteenable -> mm_interconnect_1:clock_crossing_bridge_m0_byteenable
	wire         clock_crossing_bridge_m0_readdatavalid;                    // mm_interconnect_1:clock_crossing_bridge_m0_readdatavalid -> clock_crossing_bridge:m0_readdatavalid
	wire  [31:0] clock_crossing_bridge_m0_writedata;                        // clock_crossing_bridge:m0_writedata -> mm_interconnect_1:clock_crossing_bridge_m0_writedata
	wire         clock_crossing_bridge_m0_write;                            // clock_crossing_bridge:m0_write -> mm_interconnect_1:clock_crossing_bridge_m0_write
	wire   [0:0] clock_crossing_bridge_m0_burstcount;                       // clock_crossing_bridge:m0_burstcount -> mm_interconnect_1:clock_crossing_bridge_m0_burstcount
	wire         mm_interconnect_1_ledg_s1_chipselect;                      // mm_interconnect_1:ledg_s1_chipselect -> ledg:chipselect
	wire  [31:0] mm_interconnect_1_ledg_s1_readdata;                        // ledg:readdata -> mm_interconnect_1:ledg_s1_readdata
	wire   [1:0] mm_interconnect_1_ledg_s1_address;                         // mm_interconnect_1:ledg_s1_address -> ledg:address
	wire         mm_interconnect_1_ledg_s1_write;                           // mm_interconnect_1:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_1_ledg_s1_writedata;                       // mm_interconnect_1:ledg_s1_writedata -> ledg:writedata
	wire         mm_interconnect_1_ledr_s1_chipselect;                      // mm_interconnect_1:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_1_ledr_s1_readdata;                        // ledr:readdata -> mm_interconnect_1:ledr_s1_readdata
	wire   [1:0] mm_interconnect_1_ledr_s1_address;                         // mm_interconnect_1:ledr_s1_address -> ledr:address
	wire         mm_interconnect_1_ledr_s1_write;                           // mm_interconnect_1:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_1_ledr_s1_writedata;                       // mm_interconnect_1:ledr_s1_writedata -> ledr:writedata
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                         // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [1:0] mm_interconnect_1_key_s1_address;                          // mm_interconnect_1:key_s1_address -> key:address
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                          // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                           // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_i2c_scl_s1_chipselect;                   // mm_interconnect_1:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_readdata;                     // i2c_scl:readdata -> mm_interconnect_1:i2c_scl_s1_readdata
	wire   [1:0] mm_interconnect_1_i2c_scl_s1_address;                      // mm_interconnect_1:i2c_scl_s1_address -> i2c_scl:address
	wire         mm_interconnect_1_i2c_scl_s1_write;                        // mm_interconnect_1:i2c_scl_s1_write -> i2c_scl:write_n
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_writedata;                    // mm_interconnect_1:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire         mm_interconnect_1_i2c_sda_s1_chipselect;                   // mm_interconnect_1:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_readdata;                     // i2c_sda:readdata -> mm_interconnect_1:i2c_sda_s1_readdata
	wire   [1:0] mm_interconnect_1_i2c_sda_s1_address;                      // mm_interconnect_1:i2c_sda_s1_address -> i2c_sda:address
	wire         mm_interconnect_1_i2c_sda_s1_write;                        // mm_interconnect_1:i2c_sda_s1_write -> i2c_sda:write_n
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_writedata;                    // mm_interconnect_1:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [altpll_audio:reset, altpll_sys:reset, mm_interconnect_0:altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         nios2_gen2_debug_reset_request_reset;                      // nios2_gen2:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [audio:reset, mm_interconnect_0:audio_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [clock_crossing_bridge:m0_reset, i2c_scl:reset_n, i2c_sda:reset_n, key:reset_n, ledg:reset_n, ledr:reset_n, mm_interconnect_1:clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset, sw:reset_n]
	wire         rst_controller_003_reset_out_reset;                        // rst_controller_003:reset_out -> [clock_crossing_bridge:s0_reset, data_buffer:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, onchip_memory2:reset, rst_translator:in_reset, sysid_qsys:reset_n, timer:reset_n]
	wire         rst_controller_003_reset_out_reset_req;                    // rst_controller_003:reset_req -> [data_buffer:reset_req, nios2_gen2:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]

	nios_core_altpll_audio altpll_audio (
		.clk                (clk_clk),                                            //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                     // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_audio_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_audio_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_audio_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_audio_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_audio_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_audio_c0_clk),                                //                    c0.clk
		.areset             (altpll_audio_areset_export),                         //        areset_conduit.export
		.locked             (altpll_audio_locked_export),                         //        locked_conduit.export
		.scandone           (),                                                   //           (terminated)
		.scandataout        (),                                                   //           (terminated)
		.phasedone          (),                                                   //           (terminated)
		.phasecounterselect (4'b0000),                                            //           (terminated)
		.phaseupdown        (1'b0),                                               //           (terminated)
		.phasestep          (1'b0),                                               //           (terminated)
		.scanclk            (1'b0),                                               //           (terminated)
		.scanclkena         (1'b0),                                               //           (terminated)
		.scandata           (1'b0),                                               //           (terminated)
		.configupdate       (1'b0)                                                //           (terminated)
	);

	nios_core_altpll_sys altpll_sys (
		.clk                (clk_clk),                                          //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                   // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_sys_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_sys_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_sys_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_sys_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_sys_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_sys_c0_clk),                                //                    c0.clk
		.c1                 (clk_sdram_clk),                                    //                    c1.clk
		.c2                 (clk_vga_clk),                                      //                    c2.clk
		.c3                 (altpll_sys_c3_clk),                                //                    c3.clk
		.areset             (altpll_sys_areset_export),                         //        areset_conduit.export
		.locked             (altpll_sys_locked_export),                         //        locked_conduit.export
		.scandone           (),                                                 //           (terminated)
		.scandataout        (),                                                 //           (terminated)
		.phasedone          (),                                                 //           (terminated)
		.phasecounterselect (4'b0000),                                          //           (terminated)
		.phaseupdown        (1'b0),                                             //           (terminated)
		.phasestep          (1'b0),                                             //           (terminated)
		.scanclk            (1'b0),                                             //           (terminated)
		.scanclkena         (1'b0),                                             //           (terminated)
		.scandata           (1'b0),                                             //           (terminated)
		.configupdate       (1'b0)                                              //           (terminated)
	);

	audio_if audio (
		.avalon_slave_address   (mm_interconnect_0_audio_avalon_slave_address),   // avalon_slave.address
		.avalon_slave_read      (mm_interconnect_0_audio_avalon_slave_read),      //             .read
		.avalon_slave_readdata  (mm_interconnect_0_audio_avalon_slave_readdata),  //             .readdata
		.avalon_slave_write     (mm_interconnect_0_audio_avalon_slave_write),     //             .write
		.avalon_slave_writedata (mm_interconnect_0_audio_avalon_slave_writedata), //             .writedata
		.clk                    (altpll_audio_c0_clk),                            //        clock.clk
		.reset                  (rst_controller_001_reset_out_reset),             //        reset.reset
		.BCLK                   (audio_bclk),                                     //  conduit_end.bclk
		.ADCLRC                 (audio_adclrc),                                   //             .adclrc
		.XCK                    (audio_xck),                                      //             .xck
		.ADCDAT                 (audio_adcdat),                                   //             .adcdat
		.DACLRC                 (audio_daclrc),                                   //             .daclrc
		.DACDAT                 (audio_dacdat)                                    //             .dacdat
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_bridge (
		.m0_clk           (altpll_sys_c3_clk),                                        //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                       // m0_reset.reset
		.s0_clk           (altpll_sys_c0_clk),                                        //   s0_clk.clk
		.s0_reset         (rst_controller_003_reset_out_reset),                       // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_bridge_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_bridge_m0_address),                         //         .address
		.m0_write         (clock_crossing_bridge_m0_write),                           //         .write
		.m0_read          (clock_crossing_bridge_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_bridge_m0_debugaccess)                      //         .debugaccess
	);

	nios_core_data_buffer data_buffer (
		.clk        (altpll_sys_c0_clk),                           //   clk1.clk
		.address    (mm_interconnect_0_data_buffer_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_buffer_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_buffer_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_buffer_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_buffer_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_buffer_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_buffer_s1_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_003_reset_out_reset_req),      //       .reset_req
		.freeze     (1'b0)                                         // (terminated)
	);

	nios_core_i2c_scl i2c_scl (
		.clk        (altpll_sys_c3_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_export)                           // external_connection.export
	);

	nios_core_i2c_sda i2c_sda (
		.clk        (altpll_sys_c3_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_export)                           // external_connection.export
	);

	nios_core_jtag_uart jtag_uart (
		.clk            (altpll_sys_c0_clk),                                         //               clk.clk
		.rst_n          (~rst_controller_003_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios_core_key key (
		.clk      (altpll_sys_c3_clk),                   //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_1_key_s1_address),    //                  s1.address
		.readdata (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port  (key_export)                           // external_connection.export
	);

	nios_core_ledg ledg (
		.clk        (altpll_sys_c3_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_export)                           // external_connection.export
	);

	nios_core_ledr ledr (
		.clk        (altpll_sys_c3_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	nios_core_nios2_gen2 nios2_gen2 (
		.clk                                 (altpll_sys_c0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_003_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_003_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	nios_core_onchip_memory2 onchip_memory2 (
		.clk        (altpll_sys_c0_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_003_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	nios_core_sw sw (
		.clk      (altpll_sys_c3_clk),                   //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_1_sw_s1_address),     //                  s1.address
		.readdata (mm_interconnect_1_sw_s1_readdata),    //                    .readdata
		.in_port  (sw_export)                            // external_connection.export
	);

	nios_core_sysid_qsys sysid_qsys (
		.clock    (altpll_sys_c0_clk),                                   //           clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	nios_core_timer timer (
		.clk        (altpll_sys_c0_clk),                     //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	nios_core_mm_interconnect_0 mm_interconnect_0 (
		.altpll_audio_c0_clk                                          (altpll_audio_c0_clk),                                       //                                        altpll_audio_c0.clk
		.altpll_sys_c0_clk                                            (altpll_sys_c0_clk),                                         //                                          altpll_sys_c0.clk
		.clk_50_clk_clk                                               (clk_clk),                                                   //                                             clk_50_clk.clk
		.altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // altpll_sys_inclk_interface_reset_reset_bridge_in_reset.reset
		.audio_reset_reset_bridge_in_reset_reset                      (rst_controller_001_reset_out_reset),                        //                      audio_reset_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset                 (rst_controller_003_reset_out_reset),                        //                 nios2_gen2_reset_reset_bridge_in_reset.reset
		.nios2_gen2_data_master_address                               (nios2_gen2_data_master_address),                            //                                 nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                           (nios2_gen2_data_master_waitrequest),                        //                                                       .waitrequest
		.nios2_gen2_data_master_byteenable                            (nios2_gen2_data_master_byteenable),                         //                                                       .byteenable
		.nios2_gen2_data_master_read                                  (nios2_gen2_data_master_read),                               //                                                       .read
		.nios2_gen2_data_master_readdata                              (nios2_gen2_data_master_readdata),                           //                                                       .readdata
		.nios2_gen2_data_master_readdatavalid                         (nios2_gen2_data_master_readdatavalid),                      //                                                       .readdatavalid
		.nios2_gen2_data_master_write                                 (nios2_gen2_data_master_write),                              //                                                       .write
		.nios2_gen2_data_master_writedata                             (nios2_gen2_data_master_writedata),                          //                                                       .writedata
		.nios2_gen2_data_master_debugaccess                           (nios2_gen2_data_master_debugaccess),                        //                                                       .debugaccess
		.nios2_gen2_instruction_master_address                        (nios2_gen2_instruction_master_address),                     //                          nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest                    (nios2_gen2_instruction_master_waitrequest),                 //                                                       .waitrequest
		.nios2_gen2_instruction_master_read                           (nios2_gen2_instruction_master_read),                        //                                                       .read
		.nios2_gen2_instruction_master_readdata                       (nios2_gen2_instruction_master_readdata),                    //                                                       .readdata
		.nios2_gen2_instruction_master_readdatavalid                  (nios2_gen2_instruction_master_readdatavalid),               //                                                       .readdatavalid
		.altpll_audio_pll_slave_address                               (mm_interconnect_0_altpll_audio_pll_slave_address),          //                                 altpll_audio_pll_slave.address
		.altpll_audio_pll_slave_write                                 (mm_interconnect_0_altpll_audio_pll_slave_write),            //                                                       .write
		.altpll_audio_pll_slave_read                                  (mm_interconnect_0_altpll_audio_pll_slave_read),             //                                                       .read
		.altpll_audio_pll_slave_readdata                              (mm_interconnect_0_altpll_audio_pll_slave_readdata),         //                                                       .readdata
		.altpll_audio_pll_slave_writedata                             (mm_interconnect_0_altpll_audio_pll_slave_writedata),        //                                                       .writedata
		.altpll_sys_pll_slave_address                                 (mm_interconnect_0_altpll_sys_pll_slave_address),            //                                   altpll_sys_pll_slave.address
		.altpll_sys_pll_slave_write                                   (mm_interconnect_0_altpll_sys_pll_slave_write),              //                                                       .write
		.altpll_sys_pll_slave_read                                    (mm_interconnect_0_altpll_sys_pll_slave_read),               //                                                       .read
		.altpll_sys_pll_slave_readdata                                (mm_interconnect_0_altpll_sys_pll_slave_readdata),           //                                                       .readdata
		.altpll_sys_pll_slave_writedata                               (mm_interconnect_0_altpll_sys_pll_slave_writedata),          //                                                       .writedata
		.audio_avalon_slave_address                                   (mm_interconnect_0_audio_avalon_slave_address),              //                                     audio_avalon_slave.address
		.audio_avalon_slave_write                                     (mm_interconnect_0_audio_avalon_slave_write),                //                                                       .write
		.audio_avalon_slave_read                                      (mm_interconnect_0_audio_avalon_slave_read),                 //                                                       .read
		.audio_avalon_slave_readdata                                  (mm_interconnect_0_audio_avalon_slave_readdata),             //                                                       .readdata
		.audio_avalon_slave_writedata                                 (mm_interconnect_0_audio_avalon_slave_writedata),            //                                                       .writedata
		.clock_crossing_bridge_s0_address                             (mm_interconnect_0_clock_crossing_bridge_s0_address),        //                               clock_crossing_bridge_s0.address
		.clock_crossing_bridge_s0_write                               (mm_interconnect_0_clock_crossing_bridge_s0_write),          //                                                       .write
		.clock_crossing_bridge_s0_read                                (mm_interconnect_0_clock_crossing_bridge_s0_read),           //                                                       .read
		.clock_crossing_bridge_s0_readdata                            (mm_interconnect_0_clock_crossing_bridge_s0_readdata),       //                                                       .readdata
		.clock_crossing_bridge_s0_writedata                           (mm_interconnect_0_clock_crossing_bridge_s0_writedata),      //                                                       .writedata
		.clock_crossing_bridge_s0_burstcount                          (mm_interconnect_0_clock_crossing_bridge_s0_burstcount),     //                                                       .burstcount
		.clock_crossing_bridge_s0_byteenable                          (mm_interconnect_0_clock_crossing_bridge_s0_byteenable),     //                                                       .byteenable
		.clock_crossing_bridge_s0_readdatavalid                       (mm_interconnect_0_clock_crossing_bridge_s0_readdatavalid),  //                                                       .readdatavalid
		.clock_crossing_bridge_s0_waitrequest                         (mm_interconnect_0_clock_crossing_bridge_s0_waitrequest),    //                                                       .waitrequest
		.clock_crossing_bridge_s0_debugaccess                         (mm_interconnect_0_clock_crossing_bridge_s0_debugaccess),    //                                                       .debugaccess
		.data_buffer_s1_address                                       (mm_interconnect_0_data_buffer_s1_address),                  //                                         data_buffer_s1.address
		.data_buffer_s1_write                                         (mm_interconnect_0_data_buffer_s1_write),                    //                                                       .write
		.data_buffer_s1_readdata                                      (mm_interconnect_0_data_buffer_s1_readdata),                 //                                                       .readdata
		.data_buffer_s1_writedata                                     (mm_interconnect_0_data_buffer_s1_writedata),                //                                                       .writedata
		.data_buffer_s1_byteenable                                    (mm_interconnect_0_data_buffer_s1_byteenable),               //                                                       .byteenable
		.data_buffer_s1_chipselect                                    (mm_interconnect_0_data_buffer_s1_chipselect),               //                                                       .chipselect
		.data_buffer_s1_clken                                         (mm_interconnect_0_data_buffer_s1_clken),                    //                                                       .clken
		.jtag_uart_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                       .write
		.jtag_uart_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                       .read
		.jtag_uart_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                       .chipselect
		.nios2_gen2_debug_mem_slave_address                           (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),      //                             nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                             (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),        //                                                       .write
		.nios2_gen2_debug_mem_slave_read                              (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),         //                                                       .read
		.nios2_gen2_debug_mem_slave_readdata                          (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),     //                                                       .readdata
		.nios2_gen2_debug_mem_slave_writedata                         (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),    //                                                       .writedata
		.nios2_gen2_debug_mem_slave_byteenable                        (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),   //                                                       .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),  //                                                       .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),  //                                                       .debugaccess
		.onchip_memory2_s1_address                                    (mm_interconnect_0_onchip_memory2_s1_address),               //                                      onchip_memory2_s1.address
		.onchip_memory2_s1_write                                      (mm_interconnect_0_onchip_memory2_s1_write),                 //                                                       .write
		.onchip_memory2_s1_readdata                                   (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                                       .readdata
		.onchip_memory2_s1_writedata                                  (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                                       .writedata
		.onchip_memory2_s1_byteenable                                 (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                                       .byteenable
		.onchip_memory2_s1_chipselect                                 (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                                       .chipselect
		.onchip_memory2_s1_clken                                      (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                                       .clken
		.sysid_qsys_control_slave_address                             (mm_interconnect_0_sysid_qsys_control_slave_address),        //                               sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                            (mm_interconnect_0_sysid_qsys_control_slave_readdata),       //                                                       .readdata
		.timer_s1_address                                             (mm_interconnect_0_timer_s1_address),                        //                                               timer_s1.address
		.timer_s1_write                                               (mm_interconnect_0_timer_s1_write),                          //                                                       .write
		.timer_s1_readdata                                            (mm_interconnect_0_timer_s1_readdata),                       //                                                       .readdata
		.timer_s1_writedata                                           (mm_interconnect_0_timer_s1_writedata),                      //                                                       .writedata
		.timer_s1_chipselect                                          (mm_interconnect_0_timer_s1_chipselect)                      //                                                       .chipselect
	);

	nios_core_mm_interconnect_1 mm_interconnect_1 (
		.altpll_sys_c3_clk                                          (altpll_sys_c3_clk),                       //                                        altpll_sys_c3.clk
		.clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),      // clock_crossing_bridge_m0_reset_reset_bridge_in_reset.reset
		.clock_crossing_bridge_m0_address                           (clock_crossing_bridge_m0_address),        //                             clock_crossing_bridge_m0.address
		.clock_crossing_bridge_m0_waitrequest                       (clock_crossing_bridge_m0_waitrequest),    //                                                     .waitrequest
		.clock_crossing_bridge_m0_burstcount                        (clock_crossing_bridge_m0_burstcount),     //                                                     .burstcount
		.clock_crossing_bridge_m0_byteenable                        (clock_crossing_bridge_m0_byteenable),     //                                                     .byteenable
		.clock_crossing_bridge_m0_read                              (clock_crossing_bridge_m0_read),           //                                                     .read
		.clock_crossing_bridge_m0_readdata                          (clock_crossing_bridge_m0_readdata),       //                                                     .readdata
		.clock_crossing_bridge_m0_readdatavalid                     (clock_crossing_bridge_m0_readdatavalid),  //                                                     .readdatavalid
		.clock_crossing_bridge_m0_write                             (clock_crossing_bridge_m0_write),          //                                                     .write
		.clock_crossing_bridge_m0_writedata                         (clock_crossing_bridge_m0_writedata),      //                                                     .writedata
		.clock_crossing_bridge_m0_debugaccess                       (clock_crossing_bridge_m0_debugaccess),    //                                                     .debugaccess
		.i2c_scl_s1_address                                         (mm_interconnect_1_i2c_scl_s1_address),    //                                           i2c_scl_s1.address
		.i2c_scl_s1_write                                           (mm_interconnect_1_i2c_scl_s1_write),      //                                                     .write
		.i2c_scl_s1_readdata                                        (mm_interconnect_1_i2c_scl_s1_readdata),   //                                                     .readdata
		.i2c_scl_s1_writedata                                       (mm_interconnect_1_i2c_scl_s1_writedata),  //                                                     .writedata
		.i2c_scl_s1_chipselect                                      (mm_interconnect_1_i2c_scl_s1_chipselect), //                                                     .chipselect
		.i2c_sda_s1_address                                         (mm_interconnect_1_i2c_sda_s1_address),    //                                           i2c_sda_s1.address
		.i2c_sda_s1_write                                           (mm_interconnect_1_i2c_sda_s1_write),      //                                                     .write
		.i2c_sda_s1_readdata                                        (mm_interconnect_1_i2c_sda_s1_readdata),   //                                                     .readdata
		.i2c_sda_s1_writedata                                       (mm_interconnect_1_i2c_sda_s1_writedata),  //                                                     .writedata
		.i2c_sda_s1_chipselect                                      (mm_interconnect_1_i2c_sda_s1_chipselect), //                                                     .chipselect
		.key_s1_address                                             (mm_interconnect_1_key_s1_address),        //                                               key_s1.address
		.key_s1_readdata                                            (mm_interconnect_1_key_s1_readdata),       //                                                     .readdata
		.ledg_s1_address                                            (mm_interconnect_1_ledg_s1_address),       //                                              ledg_s1.address
		.ledg_s1_write                                              (mm_interconnect_1_ledg_s1_write),         //                                                     .write
		.ledg_s1_readdata                                           (mm_interconnect_1_ledg_s1_readdata),      //                                                     .readdata
		.ledg_s1_writedata                                          (mm_interconnect_1_ledg_s1_writedata),     //                                                     .writedata
		.ledg_s1_chipselect                                         (mm_interconnect_1_ledg_s1_chipselect),    //                                                     .chipselect
		.ledr_s1_address                                            (mm_interconnect_1_ledr_s1_address),       //                                              ledr_s1.address
		.ledr_s1_write                                              (mm_interconnect_1_ledr_s1_write),         //                                                     .write
		.ledr_s1_readdata                                           (mm_interconnect_1_ledr_s1_readdata),      //                                                     .readdata
		.ledr_s1_writedata                                          (mm_interconnect_1_ledr_s1_writedata),     //                                                     .writedata
		.ledr_s1_chipselect                                         (mm_interconnect_1_ledr_s1_chipselect),    //                                                     .chipselect
		.sw_s1_address                                              (mm_interconnect_1_sw_s1_address),         //                                                sw_s1.address
		.sw_s1_readdata                                             (mm_interconnect_1_sw_s1_readdata)         //                                                     .readdata
	);

	nios_core_irq_mapper irq_mapper (
		.clk           (altpll_sys_c0_clk),                  //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_audio_c0_clk),                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_sys_c3_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (altpll_sys_c0_clk),                      //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
